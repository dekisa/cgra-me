module cgra();
    // Specifying the ports
endmodule

