module CGRA_configurator(
    input      clock,
    input      enable,
    input      sync_reset,

    output reg bitstream,
    output reg done
);

    localparam TOTAL_NUM_BITS = 844;
	reg [0:TOTAL_NUM_BITS-1] storage = {
		1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx, // block_9_3::ConstVal
		1'bx, // block_9_3::mux_out_Config
		1'bx, // block_9_3::func_Config
		1'bx,1'bx,1'bx, // block_9_3::CGAAdresPE_mux2_Config
		1'bx,1'bx,1'bx,1'bx, // block_9_3::CGAAdresPE_mux1_Config
		1'bx,1'bx,1'bx,1'bx, // block_9_3::CGAAdresPE_mux0_Config
		1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx, // block_9_2::ConstVal
		1'bx, // block_9_2::mux_out_Config
		1'bx, // block_9_2::func_Config
		1'bx,1'bx,1'bx, // block_9_2::CGAAdresPE_mux2_Config
		1'bx,1'bx,1'bx,1'bx, // block_9_2::CGAAdresPE_mux1_Config
		1'bx,1'bx,1'bx,1'bx, // block_9_2::CGAAdresPE_mux0_Config
		1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx, // block_9_1::ConstVal
		1'bx, // block_9_1::mux_out_Config
		1'bx, // block_9_1::func_Config
		1'bx,1'bx,1'bx, // block_9_1::CGAAdresPE_mux2_Config
		1'bx,1'bx,1'bx,1'bx, // block_9_1::CGAAdresPE_mux1_Config
		1'bx,1'bx,1'bx,1'bx, // block_9_1::CGAAdresPE_mux0_Config
		1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx, // block_9_0::ConstVal
		1'bx, // block_9_0::mux_out_Config
		1'bx, // block_9_0::func_Config
		1'b0,1'b0,1'b0, // block_9_0::CGAAdresPE_mux2_Config
		1'b0,1'b0,1'b0,1'b0, // block_9_0::CGAAdresPE_mux1_Config
		1'b0,1'b0,1'b0,1'b0, // block_9_0::CGAAdresPE_mux0_Config
		1'bx, // mem_port::WriteRq
		1'bx,1'bx, // mem_port::MuxData
		1'bx,1'bx, // mem_port::MuxAddr
		1'bx, // block_7_3::rf_addr_o1
		1'bx, // block_7_3::rf_addr_o0
		1'bx, // block_7_3::rf_addr_i0
		1'b0, // block_7_3::rf_WE0
		1'bx, // block_7_2::rf_addr_o1
		1'bx, // block_7_2::rf_addr_o0
		1'bx, // block_7_2::rf_addr_i0
		1'b0, // block_7_2::rf_WE0
		1'bx, // block_7_1::rf_addr_o1
		1'bx, // block_7_1::rf_addr_o0
		1'b0, // block_7_1::rf_addr_i0
		1'b1, // block_7_1::rf_WE0
		1'b1, // block_7_0::rf_addr_o1
		1'bx, // block_7_0::rf_addr_o0
		1'bx, // block_7_0::rf_addr_i0
		1'b0, // block_7_0::rf_WE0
		1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx, // block_6_3::ConstVal
		1'bx, // block_6_3::mux_out_Config
		1'bx, // block_6_3::func_Config
		1'bx,1'bx,1'bx, // block_6_3::CGAAdresPE_mux2_Config
		1'bx,1'bx,1'bx,1'bx, // block_6_3::CGAAdresPE_mux1_Config
		1'bx,1'bx,1'bx,1'bx, // block_6_3::CGAAdresPE_mux0_Config
		1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx, // block_6_2::ConstVal
		1'bx, // block_6_2::mux_out_Config
		1'bx, // block_6_2::func_Config
		1'bx,1'bx,1'bx, // block_6_2::CGAAdresPE_mux2_Config
		1'bx,1'bx,1'bx,1'bx, // block_6_2::CGAAdresPE_mux1_Config
		1'bx,1'bx,1'bx,1'bx, // block_6_2::CGAAdresPE_mux0_Config
		1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx, // block_6_1::ConstVal
		1'b0, // block_6_1::mux_out_Config
		1'bx, // block_6_1::func_Config
		1'b0,1'b0,1'b0, // block_6_1::CGAAdresPE_mux2_Config
		1'bx,1'bx,1'bx,1'bx, // block_6_1::CGAAdresPE_mux1_Config
		1'bx,1'bx,1'bx,1'bx, // block_6_1::CGAAdresPE_mux0_Config
		1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx, // block_6_0::ConstVal
		1'b1, // block_6_0::mux_out_Config
		1'b0, // block_6_0::func_Config
		1'bx,1'bx,1'bx, // block_6_0::CGAAdresPE_mux2_Config
		1'b1,1'b0,1'b0,1'b0, // block_6_0::CGAAdresPE_mux1_Config
		1'b0,1'b0,1'b0,1'b0, // block_6_0::CGAAdresPE_mux0_Config
		1'bx, // mem_port::WriteRq
		1'bx,1'bx, // mem_port::MuxData
		1'bx,1'bx, // mem_port::MuxAddr
		1'bx, // block_4_3::rf_addr_o1
		1'bx, // block_4_3::rf_addr_o0
		1'bx, // block_4_3::rf_addr_i0
		1'b0, // block_4_3::rf_WE0
		1'bx, // block_4_2::rf_addr_o1
		1'bx, // block_4_2::rf_addr_o0
		1'bx, // block_4_2::rf_addr_i0
		1'b0, // block_4_2::rf_WE0
		1'bx, // block_4_1::rf_addr_o1
		1'bx, // block_4_1::rf_addr_o0
		1'b1, // block_4_1::rf_addr_i0
		1'b1, // block_4_1::rf_WE0
		1'b1, // block_4_0::rf_addr_o1
		1'bx, // block_4_0::rf_addr_o0
		1'b1, // block_4_0::rf_addr_i0
		1'b1, // block_4_0::rf_WE0
		1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx, // block_3_3::ConstVal
		1'bx, // block_3_3::mux_out_Config
		1'bx,1'bx,1'bx,1'bx, // block_3_3::func_Config
		1'bx,1'bx,1'bx, // block_3_3::VLIWAdresPE_mux2_Config
		1'bx,1'bx,1'bx,1'bx, // block_3_3::VLIWAdresPE_mux1_Config
		1'b1,1'b1,1'b0,1'b0, // block_3_3::VLIWAdresPE_mux0_Config
		1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx, // block_3_2::ConstVal
		1'b1, // block_3_2::mux_out_Config
		1'bx,1'bx,1'bx,1'bx, // block_3_2::func_Config
		1'bx,1'bx,1'bx, // block_3_2::VLIWAdresPE_mux2_Config
		1'bx,1'bx,1'bx,1'bx, // block_3_2::VLIWAdresPE_mux1_Config
		1'bx,1'bx,1'bx,1'bx, // block_3_2::VLIWAdresPE_mux0_Config
		1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx, // block_3_1::ConstVal
		1'b1, // block_3_1::mux_out_Config
		1'bx,1'bx,1'bx,1'bx, // block_3_1::func_Config
		1'bx,1'bx,1'bx, // block_3_1::VLIWAdresPE_mux2_Config
		1'bx,1'bx,1'bx,1'bx, // block_3_1::VLIWAdresPE_mux1_Config
		1'bx,1'bx,1'bx,1'bx, // block_3_1::VLIWAdresPE_mux0_Config
		1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1, // block_3_0::ConstVal
		1'b0, // block_3_0::mux_out_Config
		1'b0,1'b0,1'b0,1'b0, // block_3_0::func_Config
		1'b0,1'b1,1'b0, // block_3_0::VLIWAdresPE_mux2_Config
		1'b0,1'b0,1'b0,1'b1, // block_3_0::VLIWAdresPE_mux1_Config
		1'b1,1'b0,1'b0,1'b1, // block_3_0::VLIWAdresPE_mux0_Config
		1'bx, // mem_port::WriteRq
		1'bx,1'bx, // mem_port::MuxData
		1'bx,1'bx, // mem_port::MuxAddr
		1'bx, // io::OEConfig
		1'bx, // io::OEConfig
		1'bx, // io::OEConfig
		1'b1, // io::OEConfig
		1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx, // block_12_3::ConstVal
		1'bx, // block_12_3::mux_out_Config
		1'bx, // block_12_3::func_Config
		1'bx,1'bx,1'bx, // block_12_3::CGAAdresPE_mux2_Config
		1'bx,1'bx,1'bx,1'bx, // block_12_3::CGAAdresPE_mux1_Config
		1'bx,1'bx,1'bx,1'bx, // block_12_3::CGAAdresPE_mux0_Config
		1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx, // block_12_2::ConstVal
		1'bx, // block_12_2::mux_out_Config
		1'bx, // block_12_2::func_Config
		1'bx,1'bx,1'bx, // block_12_2::CGAAdresPE_mux2_Config
		1'bx,1'bx,1'bx,1'bx, // block_12_2::CGAAdresPE_mux1_Config
		1'bx,1'bx,1'bx,1'bx, // block_12_2::CGAAdresPE_mux0_Config
		1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx, // block_12_1::ConstVal
		1'bx, // block_12_1::mux_out_Config
		1'bx, // block_12_1::func_Config
		1'bx,1'bx,1'bx, // block_12_1::CGAAdresPE_mux2_Config
		1'bx,1'bx,1'bx,1'bx, // block_12_1::CGAAdresPE_mux1_Config
		1'bx,1'bx,1'bx,1'bx, // block_12_1::CGAAdresPE_mux0_Config
		1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx,1'bx, // block_12_0::ConstVal
		1'b0, // block_12_0::mux_out_Config
		1'bx, // block_12_0::func_Config
		1'b0,1'b0,1'b0, // block_12_0::CGAAdresPE_mux2_Config
		1'b0,1'b0,1'b0,1'b0, // block_12_0::CGAAdresPE_mux1_Config
		1'b0,1'b0,1'b0,1'b0, // block_12_0::CGAAdresPE_mux0_Config
		1'bx, // mem_port::WriteRq
		1'bx,1'bx, // mem_port::MuxData
		1'bx,1'bx, // mem_port::MuxAddr
		1'bx, // block_10_3::rf_addr_o1
		1'bx, // block_10_3::rf_addr_o0
		1'bx, // block_10_3::rf_addr_i0
		1'b0, // block_10_3::rf_WE0
		1'bx, // block_10_2::rf_addr_o1
		1'bx, // block_10_2::rf_addr_o0
		1'bx, // block_10_2::rf_addr_i0
		1'b0, // block_10_2::rf_WE0
		1'bx, // block_10_1::rf_addr_o1
		1'bx, // block_10_1::rf_addr_o0
		1'bx, // block_10_1::rf_addr_i0
		1'b0, // block_10_1::rf_WE0
		1'bx, // block_10_0::rf_addr_o1
		1'bx, // block_10_0::rf_addr_o0
		1'bx, // block_10_0::rf_addr_i0
		1'b0, // block_10_0::rf_WE0
		1'bx,1'bx,1'bx, // block_0_0::rf_addr_o7
		1'bx,1'bx,1'bx, // block_0_0::rf_addr_o6
		1'b0,1'b0,1'b1, // block_0_0::rf_addr_o5
		1'bx,1'bx,1'bx, // block_0_0::rf_addr_o4
		1'b0,1'b0,1'b1, // block_0_0::rf_addr_o3
		1'bx,1'bx,1'bx, // block_0_0::rf_addr_o2
		1'bx,1'bx,1'bx, // block_0_0::rf_addr_o1
		1'b0,1'b0,1'b1, // block_0_0::rf_addr_o0
		1'b0,1'b0,1'b1, // block_0_0::rf_addr_i3
		1'bx,1'bx,1'bx, // block_0_0::rf_addr_i2
		1'bx,1'bx,1'bx, // block_0_0::rf_addr_i1
		1'b0,1'b0,1'b1, // block_0_0::rf_addr_i0
		1'b1, // block_0_0::rf_WE3
		1'b0, // block_0_0::rf_WE2
		1'b0, // block_0_0::rf_WE1
		1'b1 // block_0_0::rf_WE0
	};

	reg [31:0] next_pos;
	always @(posedge clock) begin
		if (sync_reset) begin
			next_pos <= 0;
			bitstream <= 1'bx;
			done <= 0;
		end else if (next_pos >= TOTAL_NUM_BITS) begin
			done <= 1;
			bitstream <= 1'bx;
		end else if (enable) begin
			bitstream <= storage[next_pos];
			next_pos <= next_pos + 1;
		end
	end
endmodule
